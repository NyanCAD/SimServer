* test
V1 1 0 DC 1 AC 1 sin(0 5 1k)
R1 1 2 1k
C2 2 0 1u
.tran 1u 2m 0
.end
